module Weight(
    input                 clk              ,
    input                 rst_n            ,
    output signed [ 15:0] o_weight_L1_0    ,
    output signed [ 15:0] o_weight_L1_1    ,
    output signed [ 15:0] o_weight_L1_2    ,
    output signed [ 15:0] o_weight_L1_3    ,
    output signed [127:0] o_weight_L2      ,
    output signed [127:0] o_weight_L3      
    );
endmodule
